module sub_module(
  input logic clock,
  input string msg
);
endmodule
