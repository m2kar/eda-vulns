module M(inout x);
endmodule
