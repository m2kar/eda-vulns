module test(input string s);
endmodule
