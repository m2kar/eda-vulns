typedef union packed { logic a; } my_union;
module Sub(input my_union x);
endmodule
