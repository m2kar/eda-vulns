module Test(inout logic c);
endmodule
