module m(input c, output real o);
always @(posedge c) o <= 0;
endmodule
