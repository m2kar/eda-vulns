module test(input string a);
endmodule
