module M(inout logic x);
endmodule
