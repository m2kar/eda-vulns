module MixedPorts(inout wire c);
endmodule
