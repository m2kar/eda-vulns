module test_module(input string a);
endmodule
