module test_module(
  input logic clk,
  output string result
);
endmodule
