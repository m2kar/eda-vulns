module t(output string s);
endmodule
