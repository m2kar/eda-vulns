module test(output string str);
endmodule
