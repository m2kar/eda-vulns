module Test(inout c);
endmodule
