module MixPorts(
  inout  wire  c
);
  assign c = 1'bz;
endmodule
