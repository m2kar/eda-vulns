module top(output string str_out);
endmodule
