module test_module(
  output string out_str
);
endmodule
