module m;
  logic [3:0] a;
  int i;
  always_comb a[i] = 1'b1;
endmodule
