module test(input string a, output int b);
endmodule
