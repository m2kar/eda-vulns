module top(input string a);
endmodule
