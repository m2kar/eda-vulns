module test_module(output string result);
endmodule
