module test_module(input string str_in);
endmodule
