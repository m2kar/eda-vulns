module e(output string o);endmodule
