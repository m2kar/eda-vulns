module test_module(output string a);
endmodule
