module M(inout logic c);
  assign c = 0;
endmodule
