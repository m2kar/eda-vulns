module M(inout d);
endmodule
