// Minimal test case for arcilator inout port crash
// Original bug: StateType cannot handle !llhd.ref<i1> from inout port
module test(inout wire c);
endmodule
