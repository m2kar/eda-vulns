module m();
  always @(*) assert (0) else $error("");
endmodule
