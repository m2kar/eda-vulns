module example(
  output string str
);
endmodule
