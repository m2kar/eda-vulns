module m(output string s);
endmodule
