module test(output string str_out);
endmodule
