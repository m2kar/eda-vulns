module Bug(inout logic c);
endmodule
