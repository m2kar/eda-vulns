module top(inout wire p);
endmodule
