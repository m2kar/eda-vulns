module top_module(output string str_out);
endmodule
