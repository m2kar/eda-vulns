module M(inout wire c);
endmodule
