module bug(inout io);
  assign io = 1'bz;
endmodule
