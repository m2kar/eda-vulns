module m(input string s);
endmodule
