typedef union packed { logic [31:0] a; } U;
module top(output U data);
endmodule
