module InoutBug(
  inout wire c
);
endmodule
