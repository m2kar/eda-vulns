module top(output string out); endmodule
