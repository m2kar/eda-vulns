module test_module(output string str_out);
endmodule
