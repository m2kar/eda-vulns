module m(
  input union packed { logic a; } u
);
endmodule
