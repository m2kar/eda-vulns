module M(inout logic c);
endmodule
