module MixPorts(
  input  logic a,
  inout  wire  c
);
  assign c = 1'b0;
endmodule
