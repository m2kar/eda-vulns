module bug(
  output string s[1:0]
);
endmodule
