module M(input string a);
endmodule
