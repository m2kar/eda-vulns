module Mod(output string str_out);
endmodule
