typedef union packed {
  logic [31:0] a;
} my_union;

module mod1(output my_union out);
endmodule
