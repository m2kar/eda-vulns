module test(output string result);
endmodule
