typedef union packed {
  logic [7:0] a;
} u_t;

module m(input u_t i);
endmodule
