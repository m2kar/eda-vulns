module Minimal(
  inout logic c
);

endmodule
