module m(inout logic x);
endmodule
